//--------------1. module----------------------//
module top_module ( input a, input b, output out );
    mod_a g0 (a, b, out);

endmodule
